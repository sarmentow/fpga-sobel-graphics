module kernel_sobel_fd();
endmodule
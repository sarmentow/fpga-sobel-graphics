module sobel_processing_unit_uc();
endmodule
module kernel_sobel_uc();
endmodule